module models

pub struct Chapter {
pub mut:
  id string
  header string
  content string
} 
